`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:26:53 01/08/2021 
// Design Name: 
// Module Name:    CPU_R 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CPU_R(clk,rst,
     PC,PC_new,Inst_code,OP,func,rs,rt,rd,
	  Write_Reg,ALU_OP,
	  RF_A,RF_B,
	  ALU_F,ZF,CF,OF,SF,PF, //
    );


endmodule
